desc_sv=Linux RAID
