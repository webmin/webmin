desc_sv=BIND DNS-server
