desc_sv=Postfixinställningar
