majordomo_cf=Fullst�ndig s�kv�g till inst�llningsfil f�r majordomo,0
program_dir=Katalog f�r majordomo-program,0
aliases_file=Aliasfil f�r sendmail-style ,3,H�mta fr�n sendmail.cf
dynamic=Anv�nda slumptal f�r listalias,1,1-Ja,0-Nej
sort_mode=Sortera mailinglistor efter,1,1-Namn,0-Ordning de skapades i
smrsh_program_dir=Katalog med sendmail-s�kerhetsprogram,3,Var som helst
