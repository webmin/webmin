named_conf=Fullständig sökväg till filen named.conf,0
named_path=Fullständig sökväg till angiven exekverbar fil,0
pid_file=Standardplacering av PID-fil,3,/var/run/named.pid
show_list=Visa domäner som,1,0-Ikoner,1-Lista
soa_style=Serienummer,1,0-Löpande nummer,1-Datumbaserade (ÅÅÅÅMMDDnn)
records_order=Visa poster ordnade,1,1-efter namn,2-efter värde,3-efter IP,0-kronologiskt
chroot=Chroot-katalog att köra BIND under,3,Standard
start_cmd=Startkommando för BIND,3,Standard
max_zones=Maximalt antal zoner att visa,0
rev_def=Förnya bakåt är,1,0-På som standard,1-Av som standard
master_ttl=Lägga till $ttl högst upp på nya zonfiler,1,1-Ja,0-Nej
named_user=Användare att starta BIND som,3,Standard
named_group=Grupp att starta BIND som,3,Standard
master_dir=Katalog för master-zonfiler,3,Standard
slave_dir=Katalog för slav/återvändszonfiler,3,Standard
support_aaaa=Stödjer DNS för IPv6-adresser,1,0-Nej,1-Ja
allow_comments=Tillåta kommentarer för poster,1,0-Nej,1-Ja
allow_wild=Tillåta jokertecken,1,0-Nej,1-Ja
