desc_sv=Webmin-användare
