raidtab=Inställningsfil för RAID,0
mdstat=Statusfil för RAID i kärnan,0
