display_max=Maximalt antal anv�ndare och grupper som ska visas,0
user_repquota_command=Kommando f�r att visa anv�ndare p� ett filsystem,0
group_repquota_command=Kommando f�r att visa grupper p� filsystem,0
user_edquota_command=Kommando f�r att �ndra en anv�ndares quota,0
group_edquota_command=Kommando f�r att �ndra en grupps quota,0
user_quota_command=Kommando f�r att kontrollera en anv�ndares quota,0
group_quota_command=Kommando f�r att kontrollera en grupps quota,0
user_copy_command=Kommando f�r att kopiera en anv�ndares quota,0
group_copy_command=Kommando f�r att kopiera en grupps quota,0
user_quotaon_command=Kommando f�r att sl� p� anv�ndares quota,0
group_quotaon_command=Kommando f�r att sl� p� gruppers quota,0
user_quotaoff_command=Kommando f�r att sl� av anv�ndares quota,0
group_quotaoff_command=Kommando f�r att sl� av gruppers quota,0
quotacheck_command=Kommando f�r att kontrollera quota,0
user_grace_command=Kommando f�r att �ndra en anv�ndares tidsintervall f�r att �verskrida quota,0
group_grace_command=Kommando f�r att �ndra en grupps tidsintervall f�r att �verskrida quota,0
