desc_sv=Postfixinst�llningar
