desc_sv=Perl-moduler
