desc_sv=PostgreSQL-databasserver
