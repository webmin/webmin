ssleay=S&#246;kv&#228;g till openssl- eller ssleay-program,0
select=Visa moduler i,1,0-Tabell,1-Rullgardinsmeny
