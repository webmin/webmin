desc_sv=Nätverkskonfigurering
