metastat_path=Fullständig sökväg till <tt>metastat</tt>,0
metadb_path=Fullständig sökväg till <tt>metadb</tt>,0
