sort_mode=Sortera tjänster och program efter,1,0-Filordning,1-Namn,2-Uppgift
inetd_conf_file=Inetd-inställningsfil,0
inetd_dir=Inetd-inställningskatalog,3,Ingen
extended_inetd=inetd-stöd,1,0-Original,1-Basstöd,2-Utökat stöd
rpc_inetd=Inetd stödjer RPCprogram,1,1-Ja,0-Nej
ipv6=Stödjer IPv6-tjänster,1,1-Ja,0-Nej
services_file=Fil för nätverkstjänster,0
rpc_file=Fil för RPC-tjänster,0
protocols_file=Fil för nätverksprotokoll,0
rpc_protocols=Underprotokoll till RPC,0
restart_command=Kommando för att starta om inetd,0
tcpd_path=Fullständig sökväg till tcpd,3
allow_file=Fullständig sökväg till tcpd allow file,3
deny_file=Fullständig sökväg till tcpd deny file,3
