desc_sv=BIND 4 DNS-server
