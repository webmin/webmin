exports_file=Exporterar fil,0
restart_command=Kommando för att starta om mountd och nfsd,0
