exports_file=Exporterar fil,0
restart_command=Kommando f�r att starta om mountd och nfsd,0
