desc_sv=Systemdokumentation
