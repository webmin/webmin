xinetd_conf=Inst&#228;llningsfil f&#246;r Xinetd,0
protocols_file=N&#228;tverksprotokollsfil,0
pid_file=S&#246;kv&#228;g till PID-fil f&#246;r Xinetd,0
start_cmd=Kommando f&#246;r att starta xinetd,0
