desc_sv=Apache Webserver
