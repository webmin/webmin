desc_sv=Startinst�llningar f�r SysV
