standard_url=URL f&#246;r standardmodul-listan&#44;3&#44;P&#229; www.webmin.com
third_url=URL f&#246;r tredje parts moduler-lista&#44;3&#44;P&#229; www.webmin.com
warn_days=Dagar f&#246;re l&#246;senord g&#229;tt ut f&#246;r att varna anv&#228;ndare&#44;0&#44;5
