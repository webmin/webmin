ftpd_path=Fullständig sökväg till wuftpd,0
ftpaccess=Fullständig sökväg till ftpaccess-fil,0
ftpconversions=Fullständig sökväg till ftpconversions-fil,0
ftpgroups=Fullständig sökväg till ftpgroups-fil,0
ftphosts=Fullständig sökväg till ftphosts-fil,0
ftpusers=Fullständig sökväg till ftpusers-fil,0
pid_file=FTP-server-PID-fil,0
