named_conf=Fullst&#228;ndig s&#246;kv&#228;g till filen named.conf,0
named_path=Fullst&#228;ndig s&#246;kv&#228;g till angiven exekverbar fil,0
pid_file=Standardplacering av PID-fil,3,/var/run/named.pid
show_list=Visa dom&#228;ner som,1,0-Ikoner,1-Lista
soa_style=Serienummer,1,0-L&#246;pande nummer,1-Datumbaserade (&#197;&#197;&#197;&#197;MMDDnn)
records_order=Visa poster ordnade,1,1-efter namn,2-efter v&#228;rde,3-efter IP,0-kronologiskt
chroot=Chroot-katalog att k&#246;ra BIND under,3,Standard
start_cmd=Startkommando f&#246;r BIND,3,Standard
max_zones=Maximalt antal zoner att visa,0
rev_def=F&#246;rnya bak&#229;t &#228;r,1,0-P&#229; som standard,1-Av som standard
master_ttl=L&#228;gga till $ttl h&#246;gst upp p&#229; nya zonfiler,1,1-Ja,0-Nej
named_user=Anv&#228;ndare att starta BIND som,3,Standard
named_group=Grupp att starta BIND som,3,Standard
master_dir=Katalog f&#246;r master-zonfiler,3,Standard
slave_dir=Katalog f&#246;r slav/&#229;terv&#228;ndszonfiler,3,Standard
support_aaaa=St&#246;djer DNS f&#246;r IPv6-adresser,1,0-Nej,1-Ja
allow_comments=Till&#229;ta kommentarer f&#246;r poster,1,0-Nej,1-Ja
allow_wild=Till&#229;ta jokertecken,1,0-Nej,1-Ja
allow_long=Till&#229;ta l&#229;nga datornamn,1,0-Nej,1-Ja
