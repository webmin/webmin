metastat_path=Fullst�ndig s�kv�g till <tt>metastat</tt>,0
metadb_path=Fullst�ndig s�kv�g till <tt>metadb</tt>,0
