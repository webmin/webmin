desc_sv=Systemloggar
