desc_sv=Webmin-anv�ndare
