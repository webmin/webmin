inittab_file=Sökväg till inittab-fil,0
