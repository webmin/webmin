exports_file=Fil med exporterade filsystem,0
restart_command=Kommando för att starta om exportserver,0
