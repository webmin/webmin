desc_sv=Listhanterare för Majordomo
