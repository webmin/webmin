desc_sv=Hjälp om Webmin
