client_conf=Konfigurationsfil f�r NIS-klient,0
nsswitch_conf=Switchfil f�r NIS-klient,0
sources=K�llor f�r nsswitch.conf,0
securenets=P�litlig n�tverksfil,3,Ingen
