exports_file=Fil med exporterade filsystem,0
restart_command=Kommando f�r att starta om exportserver,0
