smb_conf=Inst�llningsfilen f�r Samba finns h�r,0
smb_passwd=L�senordsfilen f�r Samba finns h�r,3
samba_status_program=Fullst�ndig s�kv�g till smbstatus,0
samba_password_program=Fullst�ndig s�kv�g till smbpasswd,0
samba_server=Fullst�ndig s�kv�g till smbd,0
name_server=Fullst�ndig s�kv�g till nmbd,0
swat_path=Fullst�ndig s�kv�g till swat,3,Ingen
dont_convert=Lista �ver Unix-anv�ndare som inte ska l�ggas till samba-l�senordslistan,0
sort_mode=Sortera anv�ndare och grupper efter namn,1,1-Ja,0-Nej
start_cmd=Kommando f�r att starta Samba-servrar,3,Inget
stop_cmd=Kommando f�r att stanna Samba-servrar,3,Inget
