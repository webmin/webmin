desc_sv=Konfigurations Motor
