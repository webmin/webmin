desc_sv=Användare och grupper
