desc_sv=System- och serverstatus
