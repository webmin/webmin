desc_sv=Systemtid
