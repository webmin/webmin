cron_dir=Crontab-katalog,0
cron_get_command=Kommando för att se en användares cron-jobb,0
cron_edit_command=Kommando för att ändra en användares cron-jobb,0
cron_copy_command=Kommando för att ta emot en användares cron-jobb på stdin,0
cron_delete_command=Kommando för att ta bort en användares cron-jobb,0
cron_input=Cron stödjer inmatning till cron-jobb,1,1-Ja,0-Nej
cron_allow_file=Fil med tillåtna användare,0
cron_deny_file=Fil med förbjudna användare,0
cron_deny_all=Rättigheter utan allow- eller deny-filer,1,0-Förbjud alla,1-Förbjud alla utom root,2-Tillåt alla
vixie_cron=Stödjers Vixie-Cron-tillägg,1,1-Ja,0-Nej
system_crontab=Sökväg till Vixie-Cron:s systemcrontabfil,0
cronfiles_dir=Sökväg till extra cron-filkatalog,3,Ingen
run_parts=run-parts-kommando,0
