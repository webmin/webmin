standard_url=URL för standardmodul-listan&#44;3&#44;På www.webmin.com
third_url=URL för tredje parts moduler-lista&#44;3&#44;På www.webmin.com
warn_days=Dagar före lösenord gått ut för att varna användare&#44;0&#44;5
