resolve=Sl� upp funna serveradresser,1,1-Ja,0-Nej
scan_time=V�ntetid f�r att titta efter svar,0
