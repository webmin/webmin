host=Dator att koppla upp mot,3,Automatiskt
port=Port att koppla upp mot,3,Standard
mode=Uppkopplingstyp,1,0-Telnet,1-Secure Shell (rekommenderas)
