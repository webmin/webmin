desc_sv=Schemalagda cronjobb
