inetd_conf_file=Inetd-inst�llningsfil,0
inetd_dir=Inetd-inst�llningskatalog,3,Ingen
extended_inetd=inetd-st�d,1,0-Original,1-Basst�d,2-Ut�kat st�d
show_empty=Visa tj�nster som inte har n�got program,1,1-Ja,0-Nej
rpc_inetd=Inetd st�djer RPCprogram,1,1-Ja,0-Nej
ipv6=St�djer IPv6-tj�nster,1,1-Ja,0-Nej
sort_mode=Sortera tj�nster och program efter,1,0-Filordning,1-Namn,2-Uppgift
services_file=Fil f�r n�tverkstj�nster,0
rpc_file=Fil f�r RPC-tj�nster,0
protocols_file=Fil f�r n�tverksprotokoll,0
rpc_protocols=Underprotokoll till RPC,0
restart_command=Kommando f�r att starta om inetd,0
tcpd_path=Fullst�ndig s�kv�g till tcpd,3
allow_file=Fullst�ndig s�kv�g till tcpd allow file,3
deny_file=Fullst�ndig s�kv�g till tcpd deny file,3
