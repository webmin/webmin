desc_sv=Webmin-serverindex
