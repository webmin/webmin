hosts_file=Fil med datorer och adresser,0
