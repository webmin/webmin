standard_url=URL för standardmodul-listan,3,På www.webmin.com
third_url=URL för tredje parts moduler-lista,3,På www.webmin.com
warn_days=Dagar före lösenord gått ut för att varna användare,0,5
