ftpd_path=Fullst�ndig s�kv�g till wuftpd,0
ftpaccess=Fullst�ndig s�kv�g till ftpaccess-fil,0
ftpconversions=Fullst�ndig s�kv�g till ftpconversions-fil,0
ftpgroups=Fullst�ndig s�kv�g till ftpgroups-fil,0
ftphosts=Fullst�ndig s�kv�g till ftphosts-fil,0
ftpusers=Fullst�ndig s�kv�g till ftpusers-fil,0
pid_file=FTP-server-PID-fil,0
