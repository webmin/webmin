postfix_control_command=Fullständig sökväg till Postfix-kontrollkommando,0
postfix_config_command=Fullständig sökväg till Postfix-konfigurationskommando,0
postfix_config_file=Fullständig sökväg till Postfix-konfigurationsfil,0
postfix_aliases_table_command=Fullständig sökväg till Postfix-kommando för aliasgenerering,0
postfix_newaliases_command=Fullständig sökväg till %quot;newaliases"-kommando (sendmail-kompabilitet),0
postfix_lookup_table_command=Fullständig sökväg till kommando för Postfix-uppslagstabell (`postmap'),0
