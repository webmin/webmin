xinetd_conf=Inställningsfil för Xinetd,0
protocols_file=Nätverksprotokollsfil,0
pid_file=Sökväg till PID-fil för Xinetd,0
start_cmd=Kommando för att starta xinetd,0
