desc_sv=Skrivaradministration
