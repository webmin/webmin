lilo_conf=Sökväg till LILO-inställningsfil,0
lilo_cmd=Kommando för att ta LILO-konfigurationen i drift,0
