httpd_dir=Apacheserver-rotkatalog,0
httpd_path=S&#246;kv&#228;g till exekverbar httpd-fil,0
apachectl_path=S&#246;kv&#228;g till kommando apachectl,3,Inget
start_cmd=Kommando f&#246;r att starta apache,3,Automatisk
stop_cmd=Kommando f&#246;r att stoppa apache,3,Automatisk
show_list=Visa virtuella servrar som,1,0-Ikoner,1-Lista
show_order=Sortera virtuella servrar,1,0-konfigurationsfilordning,1-servernamn,2-IP-adress
httpd_conf=S&#246;kv&#228;g till httpd.conf,3,Automatisk
srm_conf=S&#246;kv&#228;g till srm.conf,3,Automatisk
access_conf=S&#246;kv&#228;g till access.conf,3,Automatisk
mime_types=S&#246;kv&#228;g till mime.types,3,Automatisk
virt_file=L&#228;gg till virtuella servrar i filen,3,httpd.conf
