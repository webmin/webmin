desc_sv=Partitionshanterare
