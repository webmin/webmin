client_conf=Konfigurationsfil för NIS-klient,0
nsswitch_conf=Switchfil för NIS-klient,0
securenets=Pålitlig nätverksfil,3,Ingen
