ssleay=S&#246;kv&#228;g till openssl- eller ssleay-program,0
