lease=Accepterad f�rdr�jning mellan systemtid och h�rdvarutid (sekunder),0
timeserver=Standardtidserver,3,Ingen
seconds=Systemtidsformat,1,1-MMDDTTMM����.SS,0-MMDDTTMM��
zonelink=Tidszonfil,0
zonetab=Fil med tidszoner,0
zonedir=Katalog f�r tidszonfiler,0
