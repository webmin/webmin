postfix_control_command=Fullst�ndig s�kv�g till Postfix-kontrollkommando,0
postfix_config_command=Fullst�ndig s�kv�g till Postfix-konfigurationskommando,0
postfix_config_file=Fullst�ndig s�kv�g till Postfix-konfigurationsfil,0
postfix_aliases_table_command=Fullst�ndig s�kv�g till Postfix-kommando f�r aliasgenerering,0
postfix_newaliases_command=Fullst�ndig s�kv�g till %quot;newaliases&quot;-kommando (sendmail-kompabilitet),0
postfix_lookup_table_command=Fullst�ndig s�kv�g till kommando f�r Postfix-uppslagstabell (`postmap'),0
