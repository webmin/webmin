desc_sv=Squid-proxyserver
