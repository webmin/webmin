desc_sv=MySQL-databasserver
