named_boot_file=Fil f�r prim�ra inst�llningar,0
show_list=Visa dom�ner som,1,0-Ikoner,1-Lista
soa_style=Serienummer,1,0-L�pande nummer,1-Datumbaserade (����MMDDnn)
records_order=Visa poster ordnade,1,1-efter namn,0-kronologiskt
named_pid_file=Process-ID-fil,0
named_pathname=Fullst�ndig s�kv�g till <i>named</i>,0
