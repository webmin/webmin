dfstab_file=Plats för NFS-exporterade filer,0
share_all_command=Kommando för att påbörja fildelning,0
unshare_all_command=Kommando för att avsluta fildelning,0
