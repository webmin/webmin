desc_sv=Webmin-inställningar
