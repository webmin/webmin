desc_sv=Sendmail-inst�llningar
