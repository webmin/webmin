desc_sv=Schemalagda Kommandon
