passwd_file=L�senordsfil,3,Genererad
group_file=Gruppfil,0
shadow_file=Skuggl�senordsfil,3
master_file=BSD-huvudl�senordsfil,3
gshadow_file=Skuggruppfil,3
pre_command=Kommando som ska k�ras innan �ndringar g�rs,0
post_command=Kommando som ska k�ras n�r �ndringar har gjorts,0
homedir_perms=R�ttigheter f�r nya hemkataloger,0
base_uid=L�gsta UID f�r nya anv�ndare,0
base_gid=L�gsta GID f�r nya grupper,0
default_group=Standardgrupp f�r nya anv�ndare,6,Standard
display_max=Maximalt antal anv�ndare som ska visas,0
last_count=Antal tidigare inloggningar som ska visas,3,Obegr�nsat
new_user_group=Skapa ny grupp f�r nya anv�ndare,1,1-Ja,0-Nej
skip_md5=Anv�nd inte MD5-l�senord om perl-MD5-modul fattas,1,1-Ja,0-Nej
user_files=Kopiera filer till nya hemkataloger fr�n,9,40,3
display_mode=Lista med anv�ndare och grupper inneh�ller,1,2-Primary group categorised,1-Alla uppgifter,0-Endast namn
passwd_stars=D�lja l�senord i klartext?,1,1-Ja,0-Nej
delete_only=Endast ta bort filer som �gs av anv�ndaren?,1,1-Ja,0-Nej
from_files=H�mta prim�ra grupper fr�n,1,1-Fil,0-Systemanrop
alias_check=Kontrollera sendmail-alias-krockar,1,1-Ja,0-Nej
