dhcpd_conf=Konfigurationsfil för DHCP-server,0
dhcpd_path=Exekverbar fil för DHCP-server,0
pid_file=Sökväg till PID-fil för DHCP-server,0
lease_file=Lånefil för DHCP-server,0
lease_sort=Sortera lån efter,1,0-ordning i filen,1-IP-adress,2-datornamn
hostnet_list=Visa delnät och datorer som,1,0-Ikoner,1-Lista
dhcpd_nocols=ikoner i rad,0
