packages=Lista �ver CPAN-Perl-moduler,0
cpan=Grund-URL f�r CPAN-moduler,0
