index_status=Status som ska visas i listan,1,1-Aktuell status,0-Fr�n senaste schemalagda kontroll
ping_cmd=Kommando f�r att pinga en dator,3,Inget
