desc_sv=DHCP-server
