desc_sv=SSH-inloggning
