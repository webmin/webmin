inittab_file=S�kv�g till inittab-fil,0
