cron_dir=Crontab-katalog,0
cron_get_command=Kommando f�r att se en anv�ndares cron-jobb,0
cron_edit_command=Kommando f�r att �ndra en anv�ndares cron-jobb,0
cron_copy_command=Kommando f�r att ta emot en anv�ndares cron-jobb p� stdin,0
cron_delete_command=Kommando f�r att ta bort en anv�ndares cron-jobb,0
cron_input=Cron st�djer inmatning till cron-jobb,1,1-Ja,0-Nej
cron_allow_file=Fil med till�tna anv�ndare,0
cron_deny_file=Fil med f�rbjudna anv�ndare,0
cron_deny_all=R�ttigheter utan allow- eller deny-filer,1,0-F�rbjud alla,1-F�rbjud alla utom root,2-Till�t alla
vixie_cron=St�djers Vixie-Cron-till�gg,1,1-Ja,0-Nej
system_crontab=S�kv�g till Vixie-Cron:s systemcrontabfil,0
cronfiles_dir=S�kv�g till extra cron-filkatalog,3,Ingen
run_parts=run-parts-kommando,0
