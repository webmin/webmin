desc_sv=Programpaket
