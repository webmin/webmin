dhcpd_conf=Konfigurationsfil f�r DHCP-server,0
dhcpd_path=Exekverbar fil f�r DHCP-server,0
interfaces=DHCP k�r p� interface,3,Automatiskt
pid_file=S�kv�g till PID-fil f�r DHCP-server,0
lease_file=L�nefil f�r DHCP-server,0
lease_sort=Sortera l�n efter,1,0-ordning i filen,1-IP-adress,2-datornamn
hostnet_list=Visa deln�t och datorer som,1,0-Ikoner,1-Lista
dhcpd_nocols=ikoner i rad,0
