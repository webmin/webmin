index_status=Status som ska visas i listan,1,1-Aktuell status,0-Från senaste schemalagda kontroll
