desc_sv=Inställningar för start av Linux
