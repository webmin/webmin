desc_sv=Start och avstängning
