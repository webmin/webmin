pam_dir=Katalog f�r PAM-inst�llningar,0
ignore=Filer som ska ignoreras i PAM-katalogen,0
lib_dirs=Kataloger som inneh�ller PAM-bibliotek,0
mod_equiv=Utbytbara PAM-moduler,0
