lilo_conf=S�kv�g till LILO-inst�llningsfil,0
lilo_cmd=Kommando f�r att ta LILO-konfigurationen i drift,0
