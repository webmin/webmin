desc_sv=WU-FTP-server
