desc_sv=Startinställningar för SysV
