desc_sv=CD Brännare
