default_mode=Standardformat för processlista,4,last-Senast valda,tree-Processträd,user-Sorterad efter användare,size-Sorterad efter storlek,cpu-Sorterad efter CPU,search-Sökformulär,run-Utför formulär
ps_style=Format för utmatning från PS-kommandon,1,sysv-SYSV,linux-Linux,hpux-HPUX,freebsd-FreeBSD,macos-MacOS
