lease=Accepterad fördröjning mellan systemtid och hårdvarutid (sekunder),0
timeserver=Standardtidserver,3,Ingen
seconds=Systemtidsformat,1,1-MMDDTTMMÅÅÅÅ.SS,0-MMDDTTMMÅÅ
