package_system=Pakethanteringssystem,1,rpm-RPM,pkgadd-Solaris,hpux-HPUX,freebsd-FreeBSD,slackware-Slackware,debian-Debian
update_system=Automatiskt installationssystem,1,apt-Debian APT,rhn-Redhat Network,cup-Caldera CUPDATE
