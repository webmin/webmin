desc_sv=Filsystem för diskar och nätverk
