homedir_perms=Rättigheter för nya hemkataloger,0
user_files=Kopiera filer till nya hemkataloger från,9,40,3
base_uid=Lägsta UID för nya användare,0
base_gid=Lägsta GID för nya grupper,0
new_user_group=Skapa ny grupp för nya användare,1,1-Ja,0-Nej
alias_check=Kontrollera sendmail-alias-krockar,1,1-Ja,0-Nej
delete_only=Endast ta bort filer som ägs av användaren?,1,1-Ja,0-Nej
default_group=Standardgrupp för nya användare,6,Standard
display_max=Maximalt antal användare som ska visas,0
last_count=Antal tidigare inloggningar som ska visas,3,Obegränsat
display_mode=Lista med användare och grupper innehåller,1,2-Primary group categorised,1-Alla uppgifter,0-Endast namn
passwd_stars=Dölja lösenord i klartext?,1,1-Ja,0-Nej
from_files=Hämta primära grupper från,1,1-Fil,0-Systemanrop
pre_command=Kommando som ska köras innan ändringar görs,0
post_command=Kommando som ska köras när ändringar har gjorts,0
passwd_file=Lösenordsfil,3,Genererad
group_file=Gruppfil,0
shadow_file=Skugglösenordsfil,3
master_file=BSD-huvudlösenordsfil,3
gshadow_file=Skuggruppfil,3
