resolve=Slå upp funna serveradresser,1,1-Ja,0-Nej
scan_time=Väntetid för att titta efter svar,0
