desc_sv=Filsystem f�r diskar och n�tverk
