dynamic=Använda slumptal för listalias,1,1-Ja,0-Nej
sort_mode=Sortera mailinglistor efter,1,1-Namn,0-Ordning de skapades i
majordomo_cf=Fullständig sökväg till inställningsfil för majordomo,0
program_dir=Katalog för majordomo-program,0
aliases_file=Aliasfil för sendmail-style ,10,postfix-Get from Postfix,-Get from Sendmail,Other file
smrsh_program_dir=Katalog med sendmail-säkerhetsprogram,3,Var som helst
