mysqlshow=S�kv�g till mysqlshow-kommando,0
mysqladmin=S�kv�g till mysqladmin-kommando,0
mysql=S�kv�g till mysqlkommando,0
mysqldump=S�kv�g till mysqldump-kommando,0
start_cmd=Kommando f�r att starta mysql-server,0
stop_cmd=Kommando f�r att stanna mysql-server,3,Automatiskt
mysql_libs=S�kv�g till katalog f�r delade mysql-lib,3,Ingen
login=Administrat�rens inloggningsnamn,0
pass=Administrat�rens l�senord,0
perpage=Antal rader som ska visas p� en sida,0
style=Visa databaser och tabeller som,1,1-Lista,0-Ikoner
add_mode=Anv�nd vertikalt gr�nssnitt med radtill�gg,1,1-Ja,0-Nej
host=MySQL-dator att koppla upp mot,3,Localhost
sock=MySQL-socketfil,3,Standard
