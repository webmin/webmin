desc_sv=Webmin-loggning
