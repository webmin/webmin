pam_dir=Katalog för PAM-inställningar,0
ignore=Filer som ska ignoreras i PAM-katalogen,0
lib_dirs=Kataloger som innehåller PAM-bibliotek,0
mod_equiv=Utbytbara PAM-moduler,0
