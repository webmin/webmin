desc_sv=NIS-klient och -server
