syslog_conf=S�kv�g till syslog-inst�llningsfil,0
m4_conf=Syslog-inst�llningar tolkas med m4?,1,1-Ja,0-Nej
m4_path=S�kv�g till m4,0
sync=Kunna sl� av synkning efter varje meddelande?,1,1-Ja,0-Nej
pipe=St�d f�r loggning till pipor?,1,2-Till kommandon,1-Till namngivna pipor,0-Nej
pri_dir=St�d f�r avancerat prioritetsval?,1,2-FreeBSD-typ,1-Linux-typ,0-Ingen
pri_all=St�d f�r alla prioriteter?,1,1-Ja,0-Nej
tags=St�d f�r taggade sektioner?,1,1-Ja,0-Nej
pid_file=Syslog-PID-fil,3,Ingen
syslogd=S�kv�g till syslogserver,0
facilities=Resurser som st�ds,0
lines=Standardantal rader som ska visas,0
