desc_sv=Sendmail-inställningar
