desc_sv=Egna kommandon
