smb_conf=Inställningsfilen för Samba finns här,0
smb_passwd=Lösenordsfilen för Samba finns här,3
samba_status_program=Fullständig sökväg till smbstatus,0
samba_password_program=Fullständig sökväg till smbpasswd,0
samba_server=Fullständig sökväg till smbd,0
name_server=Fullständig sökväg till nmbd,0
swat_path=Fullständig sökväg till swat,3,Ingen
dont_convert=Lista över Unix-användare som inte ska läggas till samba-lösenordslistan,0
sort_mode=Sortera användare och grupper efter namn,1,1-Ja,0-Nej
start_cmd=Kommando för att starta Samba-servrar,3,Inget
stop_cmd=Kommando för att stanna Samba-servrar,3,Inget
