desc_sv=N�tverkskonfigurering
