named_boot_file=Fil för primära inställningar,0
show_list=Visa domäner som,1,0-Ikoner,1-Lista
soa_style=Serienummer,1,0-Löpande nummer,1-Datumbaserade (ÅÅÅÅMMDDnn)
records_order=Visa poster ordnade,1,1-efter namn,0-kronologiskt
named_pid_file=Process-ID-fil,0
named_pathname=Fullständig sökväg till <i>named</i>,0
