desc_sv=Webmin-inst�llningar
