default_mode=Standardformat f�r processlista,4,last-Senast valda,tree-Processtr�d,user-Sorterad efter anv�ndare,size-Sorterad efter storlek,cpu-Sorterad efter CPU,search-S�kformul�r,run-Utf�r formul�r
ps_style=Format f�r utmatning fr�n PS-kommandon,1,sysv-SYSV,linux-Linux,hpux-HPUX,freebsd-FreeBSD,macos-MacOS
