desc_sv=Hj�lp om Webmin
