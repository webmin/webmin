login=Administrat�rskonto,0
pass=Administrat�rsl�senord,0
psql=S�kv�g till psql-kommando,0
plib=S�kv�g till delade bibliotek f�r PostgreSQL,3,Beh�vs inte
basedb=PostgreSQL-databas att starta med,0
start_cmd=Kommando f�r att starta PostgreSQL,0
stop_cmd=Kommando f�r att stanna PostgreSQL,3,D�da processen
pid_file=S�kv�g till postmaster-PID-fil,0
perpage=Antal rader som ska visas per sida,0
host=PostgreSQL-dator att koppla upp mot,3,Localhost
