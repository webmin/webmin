ssleay=Sökväg till openssl- eller ssleay-program,0
