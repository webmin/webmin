dfstab_file=Plats f�r NFS-exporterade filer,0
share_all_command=Kommando f�r att p�b�rja fildelning,0
unshare_all_command=Kommando f�r att avsluta fildelning,0
