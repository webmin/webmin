raidtab=Inst�llningsfil f�r RAID,0
mdstat=Statusfil f�r RAID i k�rnan,0
