pap_file=Fil för PAP-hemligheter,0
encrypt_pass=Kryptera lösenord i filen för hemligheter,1,1-Ja,0-Nej
