packages=Lista över CPAN-Perl-moduler,0
cpan=Grund-URL för CPAN-moduler,0
