pap_file=Fil f�r PAP-hemligheter,0
encrypt_pass=Kryptera l�senord i filen f�r hemligheter,1,1-Ja,0-Nej

