desc_sv=Anv�ndare och grupper
