desc_sv=NFS-resurser
