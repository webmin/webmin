ssleay=S�kv�g till openssl- eller ssleay-program,0
select=Visa moduler i,1,0-Tabell,1-Rullgardinsmeny
