desc_sv=Listhanterare f�r Majordomo
