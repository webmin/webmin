fstab_file=Fil med filsystem som monteras vid start,0
auto_file=NFS automonterar fil,3
autofs_file=K�rnan automonterar fil,3
long_fstypes=Anv�nda l�nga filsystemtyper,1,1-Ja,0-Nej
smbclient_path=Fullst�ndig s�kv�g till <tt>smbclient</tt>,3
nmblookup_path=Fullst�ndig s�kv�g till <tt>nmblookup</tt>,3
browse_server=Server som tillhandah�ller s�klista,3,lokal
