desc_sv=Java Filhanterare
