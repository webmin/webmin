desc_sv=Inst�llningar f�r start av Linux
