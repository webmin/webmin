desc_sv=CD Br&#228;nnare
