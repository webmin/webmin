expert=Till�t individuella k�rniv�er,1,1-Ja,0-Nej
desc=Visa funktioner med beskrivningar,1,1-Ja,0-Nej
init_base=Katalog f�r k�rniv�-kataloger,0
init_dir=Katalog f�r master-init-script,0
soft_links=L�nktyp f�r k�rniv�-filer,1,0-H�rd,1-Mjuk
order_digits=Antal siffror i utf�randeordning,0
local_script=Lokalt startkommandoscript,3
reboot_command=Kommando f�r att starta om systemet,0
shutdown_command=Kommando f�r att st�nga av systemet,0
start_stop_msg=Systemet st�djer omstarts-/avst�ngningsmeddelanden,1,0-Nej,1-Ja
inittab_id=inittab-ID f�r startk�rniv�,0
daemons_dir=Katalog f�r Caldera-demoner,3,Ingen
status_check=Visa aktuell funktionsstatus,1,2-P� index- och funktionssidor,1-Endast p� funktionssidor,0-Nej
