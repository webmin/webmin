desc_sv=Fildelning med Samba
