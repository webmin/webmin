desc_sv=Start och avst�ngning
