man_cmd=Kommando f�r att visa manualsida,0
man_cmd_sect=Kommando f�r att visa manualsida ur en speciell avdelning,0
search_cmd=Kommando f�r att leta efter sidor,0
man_dir=Katalog f�r manualsidor (MANPATH),0
list_cmd=Kommando f�r att visa s�kv�g till manualsida,0
list_cmd_sect=Kommando f�r att visa s�kv�g till manualsida ur en speciell avdelning,0
man2html_path=S�kv�g till man2html,3,Anv�nd inte man2html
doc_dir=Katalog f�r paketdokumentation,3,Ingen
howto_dir=Katalog(er) f�r HOWTO-dokument,3,Ingen
kernel_dir=Katalog f�r k�rnans dokumentation,3,Ingen
kde_dir=Katalog f�r KDE-dokumentation,3,Ingen
