squid_conf=Fullst�ndig s�kv�g till inst�llningsfil f�r squid,0
squid_start=Kommando f�r att starta squid,3,Automatiskt
squid_stop=Kommando f�r att stanna squid,3,Automatiskt
squid_path=Squid-k�rfil,0
pid_file=Fullst�ndig s�kv�g till PID-fil,0
cache_dir=Fullst�ndig s�kv�g till squid-cache-katalog,0
cachemgr_path=Squid-cachemgr.cgi-k�rfil,0
log_dir=Fullst�ndig s�kv�g till squid-loggkatalog,0
calamaris=S�kv�g till logganalyseringsprogrammet calamaris,3,Inte installerat
cal_args=Argument till calamaris-kommando,0
cal_max=Maximalt antal loggrader som ska skickas till calamaris,3,Obegr�nsat
