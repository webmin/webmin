login=Administratörskonto,0
pass=Administratörslösenord,0
psql=Sökväg till psql-kommando,0
plib=Sökväg till delade bibliotek för PostgreSQL,3,Behövs inte
basedb=PostgreSQL-databas att starta med,0
start_cmd=Kommando för att starta PostgreSQL,0
stop_cmd=Kommando för att stanna PostgreSQL,3,Döda processen
pid_file=Sökväg till postmaster-PID-fil,0
perpage=Antal rader som ska visas per sida,0
host=PostgreSQL-dator att koppla upp mot,3,Localhost
