desc_sv=PAM-autentisering
