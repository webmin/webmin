desc_sv=Processhanterare
