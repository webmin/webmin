desc_sv=Backaupp Konfigurations Filer
