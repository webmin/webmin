desc_sv=Diskquota
