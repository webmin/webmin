desc_sv=NFS-exportering
