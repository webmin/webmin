browse_server=Server som tillhandahåller söklista,3,lokal
long_fstypes=Använda långa filsystemtyper,1,1-Ja,0-Nej
fstab_file=Fil med filsystem som monteras vid start,0
auto_file=NFS automonterar fil,3
autofs_file=Kärnan automonterar fil,3
smbclient_path=Fullständig sökväg till <tt>smbclient</tt>,3
nmblookup_path=Fullständig sökväg till <tt>nmblookup</tt>,3
